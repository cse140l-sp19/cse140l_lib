
//=================================
module vbuf(
input  wire reset /*synthesis syn_useioff = 0 */,          
input  wire vram_clk ,       

input  wire [7:0] data_in /* synthesis syn_force_pads=0 syn_noprune=1*/,  
input  wire data_in_rdy ,    

output wire [7:0] data_out , 
output wire data_out_rdy
) ;


parameter CYCLES_PER_BYTE = 11'd1050;
parameter BYTES_HOLD_BY_BUFFER  = 512-32;

reg [7:0] data_out_reg;
assign data_out[7:0] = data_out_reg [7:0];

reg [10:0] l_count;  
reg [8:0] r_addr, w_addr;
wire [8:0] r_addr_wire;
assign r_addr_wire [8:0] = r_addr [8:0];


//generate byte clk
//@96MHz & 921600 baud, each byte (8 + 2 stop + 1 start) need 1045.83 cycles to go through UART
always @(posedge vram_clk) begin
    if(reset) begin
        l_count <= 0;
    end
    else begin
        if(l_count == CYCLES_PER_BYTE)
            l_count <= 0;
        else 
            l_count <= l_count+1;
    end
end

//  trig_rd_h -- trig_rd_l - data_out_rdy_h .... data_out_rdy_l
wire [7:0] data_out_reg_wire;
assign data_out_rdy = l_count [10]; 

wire trig_rd;
assign trig_rd = (&l_count[9:1]) & (~l_count[10]);

wire vram_rd_clk;
assign vram_rd_clk = l_count[4];

wire vram_wr_clk;
assign vram_wr_clk = vram_clk; //l_count[3];

always @(negedge vram_rd_clk) begin
    data_out_reg[7:0] <= data_out_reg_wire[7:0];
end

always @(posedge trig_rd) begin
    if(reset)
	    r_addr <= 0;
	else
        r_addr <= r_addr + 1;
end

wire        vram_wr_en;
assign vram_wr_en = data_in_rdy & (~vram_wr_clk); // start from negative edge //vram_wr_tap;

always @(negedge vram_wr_clk) begin
    if(reset) begin
        w_addr <= 9'h000;
        //vram_wr_tap <= 0;
    end
    else begin
        if(w_addr == BYTES_HOLD_BY_BUFFER-1)
		    w_addr <= 0;
        else if(data_in_rdy)
            w_addr <= ((w_addr + 1) & 9'h0FF);
        else
            w_addr <= w_addr;
	end

end

latticeDulPortRam mem0(
.RDATA_c(data_out_reg_wire[7:0]),  //7:0
.RADDR_c(r_addr_wire[8:0]),        //8:0
.RCLK_c(vram_rd_clk),
.RCLKE_c(1'b1),
.RE_c(1'b1),

.WADDR_c(w_addr[8:0]),
.WCLK_c (vram_wr_clk),
.WCLKE_c(vram_wr_en),
.WDATA_c(data_in[7:0]),
.WE_c (vram_wr_en)
);
endmodule

//--------------------------------
module latticeDulPortRam(
output wire [7:0] RDATA_c,
input wire [8:0] RADDR_c,
input wire RCLK_c,
input wire RCLKE_c,
input wire RE_c,


input wire [8:0] WADDR_c,
input wire WCLK_c,
input wire WCLKE_c,
input wire [7:0] WDATA_c,
input wire WE_c
);

wire [7:0] RD_Dummy;
`define ICECUBE2
`ifdef ICECUBE2
SB_RAM512x8 #(
.INIT_0 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_4 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_5 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_6 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_7 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_8 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_9 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_A (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_B (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_C (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_D (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_E (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_F (256'h485b1b2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a2a0d0a)
`else
SB_RAM40_4K #(
.INIT_0 (256'h1840194509450C000C000C000C000C000C000C000C000C000CCC0CCC0CCC0CCC),
.INIT_1 (256'h084408510C000C000C000C000C000C000C000C000C000C000CCC0CCC0CCC0CCC),
.INIT_2 (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_3 (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_4 (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_5 (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_6 (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_7 (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_8 (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_9 (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_A (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_B (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_C (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_D (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_E (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.INIT_F (256'h084408510C000C000C000C000C000C000C000C000C000C000C000C000C000C00),
.READ_MODE(32'sd1),
.WRITE_MODE(32'sd1)
`endif
) ram512X8_inst (
`ifndef ICECUBE2
.MASK(16'hxxxx),
.RADDR({2'h0, RADDR_c[8:0]}),
`else
.RADDR(RADDR_c),
`endif
.RCLK(RCLK_c),
.RCLKE(RCLKE_c),
`ifndef ICECUBE2
.RDATA({RD_Dummy[7], RDATA_c[7], RD_Dummy[6], RDATA_c[6], RD_Dummy[5], RDATA_c[5], RD_Dummy[4], RDATA_c[4], 
        RD_Dummy[3], RDATA_c[3], RD_Dummy[2], RDATA_c[2], RD_Dummy[1], RDATA_c[1], RD_Dummy[0], RDATA_c[0]}),
`else
.RDATA(RDATA_c), 
`endif
.RE(RE_c),

`ifndef ICECUBE2
.WADDR({2'h0, WADDR_c[8:0]}),
`else
.WADDR(WADDR_c),
`endif
.WCLK(WCLK_c),
.WCLKE(WCLKE_c),
`ifndef ICECUBE2
.WDATA({1'hx, WDATA_c[7], 1'hx, WDATA_c[6], 1'hx, WDATA_c[5], 1'hx, WDATA_c[4], 
        1'hx, WDATA_c[3], 1'hx, WDATA_c[2], 1'hx, WDATA_c[1], 1'hx, WDATA_c[0]}),
`else
.WDATA(WDATA_c),
`endif
.WE(WE_c)
)/* synthesis syn_noprune=1 */;

/*
//0x1B [H move to home
defparam ram512x8_inst.INIT_0 =
256'h0000000000000000000000000000000000000000000000000000000000485b1b; //esc [ H
defparam ram512x8_inst.INIT_1 =
256'h0000000000000000000000000000000000000000000000000000000000000a0d;
defparam ram512x8_inst.INIT_2 =
256'h00000000000000000000000000000000000000000000002a2a2a2a2a2a000a0d;
defparam ram512x8_inst.INIT_3 =
256'h00000000000000000000000000000000000000000000002a2a2a2a2a2a000a0d;
defparam ram512x8_inst.INIT_4 =
256'h00000000000000000000000000000000000000000000002a2a00002a2a000a0d;
defparam ram512x8_inst.INIT_5 =
256'h00000000000000000000000000000000000000000000002a2a00002a2a000a0d;
defparam ram512x8_inst.INIT_6 =
256'h00000000000000000000000000000000000000000000002a2a2a2a2a2a000a0d;
defparam ram512x8_inst.INIT_7 =
256'h00000000000000000000000000000000000000000000002a2a2a2a2a2a000a0d;
defparam ram512x8_inst.INIT_8 =
256'h00000000000000000000000000000000000000000000002a2a00002a2a000a0d;
defparam ram512x8_inst.INIT_9 =
256'h00000000000000000000000000000000000000000000002a2a00002a2a000a0d;
defparam ram512x8_inst.INIT_A =
256'h00000000000000000000000000000000000000000000002a2a2a2a2a2a000a0d;
defparam ram512x8_inst.INIT_B =
256'h00000000000000000000000000000000000000000000002a2a2a2a2a2a000a0d;
defparam ram512x8_inst.INIT_C =
256'h0000000000000000000000000000000000000000000000000000000000000a0d;
defparam ram512x8_inst.INIT_D =
256'h0000000000000000000000000000000000000000000000000000000000000a0d;
defparam ram512x8_inst.INIT_E =
256'h0000000000000000000000000000000000000000000000000000000000000a0d;
defparam ram512x8_inst.INIT_F =
256'h0000000000000000000000000000000000000000000000000000000000000a0d;
*/
endmodule

